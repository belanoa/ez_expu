import fpnew_pkg::*; 

package expu_pkg;

endpackage