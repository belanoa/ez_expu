import fpnew_pkg::*; 

package expu_pkg;
    typedef enum int unsigned { BEFORE, AFTER } regs_config_t;
endpackage